assign DRAM_ADDR = 13'bxxxxxxxxxxxxx;
assign DRAM_BA = 2'bxx;
assign DRAM_CAS_N = 1;
assign DRAM_CKE = 1'bx;
assign DRAM_CLK = 1'bx;
assign DRAM_CS_N = 1;
assign DRAM_LDQM = 1'bx;
assign DRAM_RAS_N = 1;
assign DRAM_UDQM = 1'bx;
assign DRAM_WE_N = 1;

assign HEX0 = 7'bxxxxxxx;
assign HEX1 = 7'bxxxxxxx;
assign HEX2 = 7'bxxxxxxx;
assign HEX3 = 7'bxxxxxxx;
assign HEX4 = 7'bxxxxxxx;
assign HEX5 = 7'bxxxxxxx;

assign VGA_B = 8'bxxxxxxxx;
assign VGA_G = 8'bxxxxxxxx;
assign VGA_R = 8'bxxxxxxxx;
assign VGA_BLANK_N = 1;
assign VGA_CLK = 1'bx;
assign VGA_HS = 1'bx;
assign VGA_SYNC_N = 1'bx;
assign VGA_VS = 1'bx;

assign ADC_DIN = 1'bx;
assign ADC_SCLK = 1'bx;

assign AUD_DACDAT = 1'bx;
assign AUD_XCK = 1'bx;

assign FAN_CTRL = 1'bx;

assign FPGA_I2C_SCLK = 1'bx;

assign HPS_FLASH_DCLK = 1'bx;
assign HPS_FLASH_NCSO = 1;
assign HPS_SPIM_CLK = 1'bx;
assign HPS_SPIM_MOSI = 1'bx;

assign IRDA_TXD = 1'bx;
assign TD_RESET_N = 0;
